library verilog;
use verilog.vl_types.all;
entity sam_test is
end sam_test;

library verilog;
use verilog.vl_types.all;
entity ma_test is
end ma_test;
